package tb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import agent_pkg::*;
  `include "mem_scoreboard.sv"
  `include "mem_env.sv"
  `include "mem_basic_test.sv"
endpackage